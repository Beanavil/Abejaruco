`default_nettype none

module abejaruco(input a, input b, output y);
    //
endmodule