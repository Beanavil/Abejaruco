// GNU General Public License
//
// Copyright : (c) 2023 Javier Beiro Piñón
// : (c) 2023 Beatriz Navidad Vilches
// : (c) 2023 Stefano Petrilli
//
// This file is part of Abejaruco <https:// github.com/Beanavil/Abejaruco>.
//
// Abejaruco is free software: you can redistribute it and/or modify it under
// the terms of the GNU General Public License as published by the Free
// Software Foundation, either version 3 of the License, or (at your option)
// any later version.
//
// Abejaruco is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS
// FOR A PARTICULAR PURPOSE. See the GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with Abejaruco placed on the LICENSE.md file of the root folder.
// If not, see <https:// www.gnu.org/licenses/>.

`ifndef TAG_COMPARATOR_V
`define TAG_COMPARATOR_V

module tag_comparator(
    input wire [TAG_WIDTH-1:0] input_tag,
    input wire [TAG_WIDTH-1:0] stored_tag,
    input wire valid,
    output wire hit
  );
`include "src/parameters.v"

  assign hit = valid ? (input_tag == stored_tag) : 1'b0;
endmodule

`endif
