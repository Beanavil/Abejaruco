`default_nettype none

module Abejaruco_tb(input a,
                   input b,
                   output y);
  //
endmodule
